module pc_mais_4
(pc,pc_mais_4);
input [31:0] pc;
output wire [31:0] pc_mais_4;

assign pc_mais_4 = pc + 32'd4;

endmodule
