module ADD
(ent1,ent2,saida);
input [31:0] ent1, ent2;
output wire [31:0] saida;
assign saida = ent1 + ent2;
endmodule
