library verilog;
use verilog.vl_types.all;
entity ProcessadorMips_vlg_vec_tst is
end ProcessadorMips_vlg_vec_tst;
